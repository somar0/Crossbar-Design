library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg.all;
 
entity threshold_rom is
port(	
    Clk           : in std_logic;
	Reset         : in std_logic;	
	add	          : in std_logic_vector(7 downto 0);    -- Adress
	Threshold_out : out std_logic_vector(31 downto 0)   -- Threshold Rom Output
);
end threshold_rom;



architecture rtl of threshold_rom is
    -- The Values of the Threshold Matrix
    constant Content: threshold_array(0 to alpha-1) := (
        0   => "00000000000000000000000000110110",
        1   => "00000000000000000000000100010001",
        2   => "00000000000000000000000110100101",
        3   => "00000000000000000000000110001011",
        4   => "00000000000000000000000000100010",
        5   => "00000000000000000000000100101000",
        6   => "00000000000000000000000011000110",
        7   => "00000000000000000000000100010110",
        8   => "00000000000000000000000011101111",
        9   => "00000000000000000000000101001001",
        10  => "00000000000000000000001000011110",
        11  => "00000000000000000000000001000101",
        12  => "00000000000000000000000011010011",
        13  => "00000000000000000000000000010101",
        14  => "00000000000000000000000000000110",
        15  => "00000000000000000000000111000100",
        16  => "00000000000000000000000101011111",
        17  => "00000000000000000000000010110011",
        18  => "00000000000000000000000100011000",
        19  => "00000000000000000000000001101111",
        20  => "00000000000000000000000001010110",
        21  => "00000000000000000000000111001100",
        22  => "00000000000000000000000100101101",
        23  => "00000000000000000000000101111011",
        24  => "00000000000000000000000010010000",
        25  => "00000000000000000000001000111111",
        26  => "00000000000000000000000101110111",
        27  => "00000000000000000000000110110001",
        28  => "00000000000000000000000100001001",
        29  => "00000000000000000000001000010001",
        30  => "00000000000000000000000001010100",
        31  => "00000000000000000000000100010010",
        32  => "00000000000000000000000000000110",
        33  => "00000000000000000000000010011101",
        34  => "00000000000000000000001000110111",
        35  => "00000000000000000000000001000110",
        36  => "00000000000000000000000011111100",
        37  => "00000000000000000000000010100110",
        38  => "00000000000000000000001000000101",
        39  => "00000000000000000000001000011011",
        40  => "00000000000000000000000010000111",
        41  => "00000000000000000000000101000111",
        42  => "00000000000000000000000101111110",
        43  => "00000000000000000000000111011010",
        44  => "00000000000000000000000110010001",
        45  => "00000000000000000000000001111100",
        46  => "00000000000000000000000000110100",
        47  => "00000000000000000000000000111111",
        48  => "00000000000000000000000001100100",
        49  => "00000000000000000000000111111111",
        50  => "00000000000000000000000011001000",
        51  => "00000000000000000000000011100000",
        52  => "00000000000000000000000101101011",
        53  => "00000000000000000000000101110001",
        54  => "00000000000000000000000101111110",
        55  => "00000000000000000000000000001011",
        56  => "00000000000000000000000011010001",
        57  => "00000000000000000000000000111000",
        58  => "00000000000000000000000010010010",
        59  => "00000000000000000000000010010001",
        60  => "00000000000000000000000011100000",
        61  => "00000000000000000000000011101001",
        62  => "00000000000000000000000111111100",
        63  => "00000000000000000000000000111011"
    );       
    
begin
    -- Read Process
    process(clk, Reset)
    begin
        if rising_edge(clk) then
            if( Reset = '1' ) then
                Threshold_out  <= (others => '0');
            else 
                Threshold_out  <= Content(to_integer(unsigned(add)));
            end if;
        end if;
    end process;
end rtl;

